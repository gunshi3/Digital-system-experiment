-- Copyright (C) 1991-2009 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.0 Build 184 04/29/2009 Service Pack 1 SJ Web Edition
-- Created on Mon Apr 26 11:35:28 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY exp_detect3 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        din : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC
    );
END exp_detect3;

ARCHITECTURE BEHAVIOR OF exp_detect3 IS
    TYPE type_fstate IS (s0,s1,s2,s3,s4,s5,s6);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='1') THEN
            fstate <= s0;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,din)
    BEGIN
        z <= '0';
        CASE fstate IS
            WHEN s0 =>
                IF (NOT((din = '1'))) THEN
                    reg_fstate <= s0;
                ELSIF ((din = '1')) THEN
                    reg_fstate <= s1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s0;
                END IF;
            WHEN s1 =>
                IF ((din = '1')) THEN
                    reg_fstate <= s2;
                ELSIF (NOT((din = '1'))) THEN
                    reg_fstate <= s0;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s1;
                END IF;
            WHEN s2 =>
                IF (NOT((din = '1'))) THEN
                    reg_fstate <= s0;
                ELSIF ((din = '1')) THEN
                    reg_fstate <= s3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s2;
                END IF;
            WHEN s3 =>
                IF (NOT((din = '1'))) THEN
                    reg_fstate <= s4;
                ELSIF ((din = '1')) THEN
                    reg_fstate <= s3;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s3;
                END IF;
            WHEN s4 =>
                IF (NOT((din = '1'))) THEN
                    reg_fstate <= s5;
                ELSIF ((din = '1')) THEN
                    reg_fstate <= s1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s4;
                END IF;
            WHEN s5 =>
                IF (NOT((din = '1'))) THEN
                    reg_fstate <= s0;
                ELSIF ((din = '1')) THEN
                    reg_fstate <= s6;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s5;
                END IF;
            WHEN s6 =>
                IF (NOT((din = '1'))) THEN
                    reg_fstate <= s0;
                ELSIF ((din = '1')) THEN
                    reg_fstate <= s2;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= s6;
                END IF;

                IF (NOT((din = '1'))) THEN
                    z <= '1';
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    z <= '0';
                END IF;
            WHEN OTHERS => 
                z <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
